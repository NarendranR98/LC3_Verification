package decode_out_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "src/decode_out_configuration.sv" 
    `include "src/decode_out_transaction.sv" 
    `include "src/decode_out_monitor.sv"
    `include "src/decode_out_agent.sv"
endpackage