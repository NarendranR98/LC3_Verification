package decode_test_pkg;
 import uvm_pkg::*;
 import decode_in_pkg::*;
 `include "uvm_macros.svh"
 `include "src/test_top.sv"
endpackage