interface decode_in_if(input clock,input reset);
logic enable_decode;
logic [15:0] Instr_dout;
logic [15:0] npc_in;
endinterface